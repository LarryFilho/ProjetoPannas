LIBRARY ieee;
USE ieee.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.ALL;

PACKAGE conexao IS
	SUBTYPE reg16 IS std_logic_vector(15 downto 0);
END conexao;